`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Tsinghua University
// Engineer: Timothy-LiuXuefeng
// 
// Create Date: 2021/07/08 12:16:51
// Design Name: PipelineCPU
// Module Name: PipelineCPU
// Project Name: PipelineCPU
// Target Devices: xc7a35tcpg236-1
// Tool Versions: Vivado 2017.3
// Description: Top design module.
// 
// Dependencies: None
// 
// Revision: None
// Revision 0.01 - File Created
// Additional Comments: None
// 
//////////////////////////////////////////////////////////////////////////////////


module PipelineCPU
(
    input wire clk,
    input wire reset,
    output wire [7:0] leds,
    output wire [3:0] AN,
    output wire [3:0] BCD
);

endmodule
